module four_input_and_gate(input A, B, C, D, output E);

    assign E = A & B & C & D;        
endmodule