module four_input_and(input A, B, C, D, output out_and);

    assign out_and = A & B & C & D;

endmodule